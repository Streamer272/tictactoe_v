module content

pub const (
	covered = `■`
	x = `X`
	y = `Y`
)
