module field

pub enum Direction {
	up
	down
	left
	right
}
