module main

import field { new_field }

fn main() {
	field := new_field()
	println("Field: $field")
}
