module box

pub enum Content {
	empty
	x
	y
}
