module content

pub enum Content {
	covered
	selected
	uncovered_x
	uncovered_o
}
