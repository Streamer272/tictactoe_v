module direction

pub enum Direction {
	up
	down
	left
	right
}
